module testbench(
    clk

    );
    
    
    
    
    
    
    
    
endmodule

module testbench(
    clk

    );
    
    
    
    
    
    
    
    
endmodule